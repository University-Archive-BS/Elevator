`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AUT-CEIT
// Engineer: Ali Nazari
// Create Date:    16:23:13 01/21/2019 
// Module Name:    elevator 
// Project Name: Smart-Elevator 
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module elevator(
    );


endmodule
